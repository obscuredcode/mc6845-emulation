module hex_segment(in)

input reg[0:3] in;

always
begin
	
end

endmodule