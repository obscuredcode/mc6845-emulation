module hex_segment(input in);

//input reg[0:3] in;

always
begin
	
end

endmodule